library verilog;
use verilog.vl_types.all;
entity chip_top is
end chip_top;
